module alu_plus(input [9:0] a, b , output [9:0]out);
  assign out = a + b;
endmodule
library verilog;
use verilog.vl_types.all;
entity memory is
    port(
        clk             : in     vl_logic;
        adr             : in     vl_logic_vector(9 downto 0);
        \out\           : out    vl_logic_vector(15 downto 0);
        write_data      : in     vl_logic_vector(15 downto 0);
        mem_read        : in     vl_logic;
        mem_write       : in     vl_logic
    );
end memory;
